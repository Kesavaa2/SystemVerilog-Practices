interface inter;

  logic clk,data,reset,q;
  
endinterface
