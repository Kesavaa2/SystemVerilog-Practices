interface operation;
  
  logic a,b,c;
  
  bit sum,carry;

endinterface
  
