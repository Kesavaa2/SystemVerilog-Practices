interface dff_intf;

  logic clk;
  logic rst;
  logic d;
  logic q;
  
endinterface
