interface intf;
  logic a,b,c,sum,Cout;
endinterface
