class transaction;

  rand bit data;
  bit reset;
  bit q;

endclass
